-- Simple interface to tx side of transactor...
-- Even simpler, but now multi-buffer RAM!
--
-- Dave Sankey, September 2012

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity udp_txtransactor_if is
  generic(
    BUFWIDTH: natural := 0
  );
  port (
    mac_clk: in std_logic;
    rst_macclk: in std_logic;
--
    pkt_resend: in std_logic;
    resend_pkt_id: in std_logic_vector(15 downto 0);
--
    ipbus_out_hdr: in std_logic_vector(31 downto 0);
    ipbus_out_valid: in std_logic;
    tx_read_buffer: in std_logic_vector(BUFWIDTH - 1 downto 0);
--
    udpram_busy: in std_logic;
    clean_buf: in std_logic_vector(2**BUFWIDTH - 1 downto 0);
--
    req_resend: out std_logic;
    resend_buf: out std_logic_vector(BUFWIDTH - 1 downto 0);
    udpram_sent: out std_logic
  );
end udp_txtransactor_if;

architecture simple of udp_txtransactor_if is

  type pktid_buf is array (2**BUFWIDTH - 1 downto 0) of std_logic_vector(15 downto 0);
  signal pkt_id_buf: pktid_buf;

begin

pkt_id_block: process (mac_clk)
  begin
    if rising_edge(mac_clk) then
      if rst_macclk = '1' then
	pkt_id_buf <= (Others => (Others => '0'));
      elsif ipbus_out_valid = '1' then
	pkt_id_buf(to_integer(unsigned(tx_read_buffer))) <= ipbus_out_hdr(23 downto 8);
      end if;
    end if;
  end process;

resend_block: process (mac_clk)
  variable req_resend_i: std_logic;
  variable resend_buf_i: std_logic_vector(BUFWIDTH - 1 downto 0);
  begin
    if rising_edge(mac_clk) then
      req_resend_i := '0';
      resend_buf_i := (Others => '0');
      if pkt_resend = '1' then
        for i in 0 to 2**BUFWIDTH - 1 loop
          if pkt_id_buf(i) = resend_pkt_id and clean_buf(i) = '1' then
	    req_resend_i := '1';
	    resend_buf_i := std_logic_vector(to_unsigned(i, BUFWIDTH));
	  end if;
        end loop;
      end if;
      req_resend <= req_resend_i
-- pragma translate_off
      after 4 ns
-- pragma translate_on
      ;
      resend_buf <= resend_buf_i
-- pragma translate_off
      after 4 ns
-- pragma translate_on
      ;
    end if;
  end process;

sent_block: process (mac_clk)
  variable last_busy: std_logic;
  begin
    if rising_edge(mac_clk) then
      udpram_sent <= last_busy and not udpram_busy
-- pragma translate_off
      after 4 ns
-- pragma translate_on
      ;
      last_busy := udpram_busy;
    end if;
  end process;

end simple;
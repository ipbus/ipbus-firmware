---------------------------------------------------------------------------------
--
--   Copyright 2017 - Rutherford Appleton Laboratory and University of Bristol
--
--   Licensed under the Apache License, Version 2.0 (the "License");
--   you may not use this file except in compliance with the License.
--   You may obtain a copy of the License at
--
--       http://www.apache.org/licenses/LICENSE-2.0
--
--   Unless required by applicable law or agreed to in writing, software
--   distributed under the License is distributed on an "AS IS" BASIS,
--   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--   See the License for the specific language governing permissions and
--   limitations under the License.
--
--                                     - - -
--
--   Additional information about ipbus-firmare and the list of ipbus-firmware
--   contacts are available at
--
--       https://ipbus.web.cern.ch/ipbus
--
---------------------------------------------------------------------------------


-- eth_7s_1000basex_gtp
--
-- Contains the instantiation of the Xilinx MAC & 1000baseX pcs/pma & GTP transceiver cores
--
-- This version is for the artix GTP transceivers, and has the GTPE2_COMMON included in this block.
-- Various PLL clock outputs are therefore provided for use by other MGTs in the same quad.
--
-- Do not change signal names in here without corresponding alteration to the timing contraints file
--
-- Dave Newbold, January 2016

library ieee;
use ieee.std_logic_1164.all;

library unisim;
use unisim.VComponents.all;

entity bp_eth_7s_1000basex_gtp_shared_logic_in is
	port(
		gt_txp, gt_txn: out std_logic;
		gt_rxp, gt_rxn: in std_logic;

		tx_data: in std_logic_vector(7 downto 0);
		tx_valid: in std_logic;
		tx_last: in std_logic;
		tx_error: in std_logic;
		tx_ready: out std_logic;
		rx_data: out std_logic_vector(7 downto 0);
		rx_valid: out std_logic;
		rx_last: out std_logic;
		rx_error: out std_logic;
		
        -- Replacing clk_iface record structure.
        clk125          : in std_logic;
        clk125_fr      : in std_logic;
        rst_eth         : in std_logic;
        clk_indep       : in std_logic;
        
        -- Replacing phy_iface record structure.
        pma_reset               : in std_logic;
        gt0_pll0outclk_in       : in std_logic;
        gt0_pll0outrefclk_in    : in std_logic;
        gt0_pll1outclk_in       : in std_logic;
        gt0_pll1outrefclk_in    : in std_logic;
        gt0_pll0lock_in         : in std_logic;
        gt0_pll0refclklost_in   : in std_logic;
        user_clk                : in std_logic;
        gtrefclk                : in std_logic;
        mmcm_locked             : in std_logic;
        locked                  : out std_logic
	);

end bp_eth_7s_1000basex_gtp_shared_logic_in;

architecture rtl of bp_eth_7s_1000basex_gtp_shared_logic_in is

	COMPONENT temac_gbe_v9_0
		PORT (
			gtx_clk : IN STD_LOGIC;
			glbl_rstn : IN STD_LOGIC;
			rx_axi_rstn : IN STD_LOGIC;
			tx_axi_rstn : IN STD_LOGIC;
			rx_statistics_vector : OUT STD_LOGIC_VECTOR(27 DOWNTO 0);
			rx_statistics_valid : OUT STD_LOGIC;
			rx_mac_aclk : OUT STD_LOGIC;
			rx_reset : OUT STD_LOGIC;
			rx_axis_mac_tdata : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			rx_axis_mac_tvalid : OUT STD_LOGIC;
			rx_axis_mac_tlast : OUT STD_LOGIC;
			rx_axis_mac_tuser : OUT STD_LOGIC;
			tx_ifg_delay : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			tx_statistics_vector : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			tx_statistics_valid : OUT STD_LOGIC;
			tx_mac_aclk : OUT STD_LOGIC;
			tx_reset : OUT STD_LOGIC;
			tx_axis_mac_tdata : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			tx_axis_mac_tvalid : IN STD_LOGIC;
			tx_axis_mac_tlast : IN STD_LOGIC;
			tx_axis_mac_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
			tx_axis_mac_tready : OUT STD_LOGIC;
			pause_req : IN STD_LOGIC;
			pause_val : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			speedis100 : OUT STD_LOGIC;
			speedis10100 : OUT STD_LOGIC;
			gmii_txd : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			gmii_tx_en : OUT STD_LOGIC;
			gmii_tx_er : OUT STD_LOGIC;
			gmii_rxd : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			gmii_rx_dv : IN STD_LOGIC;
			gmii_rx_er : IN STD_LOGIC;
			rx_configuration_vector : IN STD_LOGIC_VECTOR(79 DOWNTO 0);
			tx_configuration_vector : IN STD_LOGIC_VECTOR(79 DOWNTO 0)
		);
	END COMPONENT;

	signal gmii_txd, gmii_rxd: std_logic_vector(7 downto 0);
	signal gmii_tx_en, gmii_tx_er, gmii_rx_dv, gmii_rx_er: std_logic;
	signal rx_rec_clk, rx_rec_clk_i: std_logic;
	signal rstn, phy_done, locked_int: std_logic;
	
	attribute mark_debug: string;
    attribute mark_debug of rstn, locked_int, mmcm_locked, phy_done: signal is "True";
    attribute mark_debug of gmii_txd, gmii_tx_en, gmii_tx_er, gmii_rxd, gmii_rx_dv, gmii_rx_er : signal is "True";
	
begin

	process(clk125)
	begin
		if rising_edge(clk125) then
			locked_int <= mmcm_locked and phy_done;
		end if;
	end process;

    locked <= locked_int;
	rstn <= not (not locked_int or rst_eth);

	mac: temac_gbe_v9_0
		port map(
			gtx_clk => clk125,
			glbl_rstn => rstn,
			rx_axi_rstn => '1',
			tx_axi_rstn => '1',
			rx_statistics_vector => open,
			rx_statistics_valid => open,
			rx_mac_aclk => open,
			rx_reset => open,
			rx_axis_mac_tdata => rx_data,
			rx_axis_mac_tvalid => rx_valid,
			rx_axis_mac_tlast => rx_last,
			rx_axis_mac_tuser => rx_error,
			tx_ifg_delay => X"00",
			tx_statistics_vector => open,
			tx_statistics_valid => open,
			tx_mac_aclk => open,
			tx_reset => open,
			tx_axis_mac_tdata => tx_data,
			tx_axis_mac_tvalid => tx_valid,
			tx_axis_mac_tlast => tx_last,
			tx_axis_mac_tuser(0) => tx_error,
			tx_axis_mac_tready => tx_ready,
			pause_req => '0',
			pause_val => X"0000",
			gmii_txd => gmii_txd,
			gmii_tx_en => gmii_tx_en,
			gmii_tx_er => gmii_tx_er,
			gmii_rxd => gmii_rxd,
			gmii_rx_dv => gmii_rx_dv,
			gmii_rx_er => gmii_rx_er,
			rx_configuration_vector => X"0000_0000_0000_0000_0812",
			tx_configuration_vector => X"0000_0000_0000_0000_0012"
		);

    bp_phy : entity work.gig_eth_pcs_pma_basex_gtp_no_shared_logic
        port map(
            gtrefclk_bufg => clk125_fr,
            gtrefclk => gtrefclk,
            
            txp => gt_txp,
            txn => gt_txn,
            rxp => gt_rxp,
            rxn => gt_rxn,
            
            resetdone => phy_done,
            cplllock => open,
            
            mmcm_reset => open,
            
            txoutclk => open,
            rxoutclk => rx_rec_clk,
            
            userclk => user_clk,
            userclk2 => clk125,
            
            rxuserclk => rx_rec_clk_i,
            rxuserclk2 => rx_rec_clk_i,
            
            independent_clock_bufg => clk_indep,
            pma_reset => pma_reset,
            mmcm_locked => mmcm_locked,
            
            gmii_txd => gmii_txd,
            gmii_tx_en => gmii_tx_en,
            gmii_tx_er => gmii_tx_er,
            gmii_rxd => gmii_rxd,
            gmii_rx_dv => gmii_rx_dv,
            gmii_rx_er => gmii_rx_er,
            gmii_isolate => open,
            
            configuration_vector => "00000",
            status_vector => open,
            reset => rst_eth,
            
            signal_detect => '1',
            
            gt0_pll0outclk_in => gt0_pll0outclk_in,
            gt0_pll0outrefclk_in => gt0_pll0outrefclk_in,
            gt0_pll1outclk_in => gt0_pll1outclk_in,
            gt0_pll1outrefclk_in => gt0_pll1outrefclk_in,
            gt0_pll0lock_in => gt0_pll0lock_in,
            gt0_pll0refclklost_in => gt0_pll0refclklost_in,
            gt0_pll0reset_out => open
        );
        
        -- Clocks
        bufg_rx_clk: BUFG
        port map(
            i =>  rx_rec_clk,
            o =>  rx_rec_clk_i
        );
end rtl;

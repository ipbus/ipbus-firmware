-------------------------------------------------------------------------------
--   __  __ 
--  /   /\/   / 
-- /__/  \   /    Vendor: Xilinx 
-- \   \   \/     Version : 1.2
--  \   \         Application : RocketIO GTX Wizard 
--  /   /         Filename : rocketio_wrapper_gtx_vhdl_tile.vhd
-- /__/   /\      Timestamp : 02/08/2005 09:12:43
-- \   \  /  \ 
--  \__\/\__\ 
--
--
-- Module ROCKETIO_WRAPPER_GTX_TILE (a GTX Tile Wrapper)
-- Generated by Xilinx RocketIO GTX Wizard

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***************************** Entity Declaration ****************************

entity ROCKETIO_WRAPPER_GTX_TILE is
generic
(
    -- Simulation attributes
    TILE_SIM_GTXRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    TILE_SIM_PLL_PERDIV2         : bit_vector:= x"0c8"; -- Set to the VCO Unit Interval time 

    -- Channel bonding attributes
    TILE_CHAN_BOND_MODE_0        : string    := "OFF";  -- "MASTER", "SLAVE", or "OFF"
    TILE_CHAN_BOND_LEVEL_0       : integer   := 0;     -- 0 to 7. See UG for details
    
    TILE_CHAN_BOND_MODE_1        : string    := "OFF";  -- "MASTER", "SLAVE", or "OFF"
    TILE_CHAN_BOND_LEVEL_1       : integer   := 0      -- 0 to 7. See UG for details
);
port 
(
    ------------------------ Loopback and Powerdown Ports ----------------------
    LOOPBACK0_IN                            : in   std_logic_vector(2 downto 0);
    LOOPBACK1_IN                            : in   std_logic_vector(2 downto 0);
    RXPOWERDOWN0_IN                         : in   std_logic_vector(1 downto 0);
    TXPOWERDOWN0_IN                         : in   std_logic_vector(1 downto 0);
    RXPOWERDOWN1_IN                         : in   std_logic_vector(1 downto 0);    
    TXPOWERDOWN1_IN                         : in   std_logic_vector(1 downto 0);    
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    RXCHARISCOMMA0_OUT                      : out  std_logic;
    RXCHARISK0_OUT                          : out  std_logic;
    RXDISPERR0_OUT                          : out  std_logic;
    RXNOTINTABLE0_OUT                       : out  std_logic;
    RXRUNDISP0_OUT                          : out  std_logic;
    RXCHARISCOMMA1_OUT                      : out  std_logic;
    RXCHARISK1_OUT                          : out  std_logic;
    RXDISPERR1_OUT                          : out  std_logic;
    RXNOTINTABLE1_OUT                       : out  std_logic;
    RXRUNDISP1_OUT                          : out  std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    RXCLKCORCNT0_OUT                        : out  std_logic_vector(2 downto 0);
    RXCLKCORCNT1_OUT                        : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    RXENMCOMMAALIGN0_IN                     : in   std_logic;
    RXENMCOMMAALIGN1_IN                     : in   std_logic;
    RXENPCOMMAALIGN0_IN                     : in   std_logic;
    RXENPCOMMAALIGN1_IN                     : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    RXDATA0_OUT                             : out  std_logic_vector(7 downto 0);
    RXDATA1_OUT                             : out  std_logic_vector(7 downto 0);
    RXRECCLK0_OUT                           : out  std_logic;
    RXRECCLK1_OUT                           : out  std_logic;
    RXRESET0_IN                             : in   std_logic;
    RXRESET1_IN                             : in   std_logic;
    RXUSRCLK0_IN                            : in   std_logic;
    RXUSRCLK1_IN                            : in   std_logic;
    RXUSRCLK20_IN                           : in   std_logic;
    RXUSRCLK21_IN                           : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    RXELECIDLE0_OUT                         : out  std_logic;
    RXELECIDLE1_OUT                         : out  std_logic;
    RXN0_IN                                 : in   std_logic;
    RXN1_IN                                 : in   std_logic;
    RXP0_IN                                 : in   std_logic;
    RXP1_IN                                 : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    RXBUFRESET0_IN                          : in   std_logic;
    RXBUFRESET1_IN                          : in   std_logic;
    RXBUFSTATUS0_OUT                        : out  std_logic_vector(2 downto 0);
    RXBUFSTATUS1_OUT                        : out  std_logic_vector(2 downto 0);
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    CLKIN_IN                                : in   std_logic;
    GTXRESET_IN                             : in   std_logic;
    PLLLKDET_OUT                            : out  std_logic;
    REFCLKOUT_OUT                           : out  std_logic;
    RESETDONE0_OUT                          : out  std_logic;
    RESETDONE1_OUT                          : out  std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TXCHARDISPMODE0_IN                      : in   std_logic;
    TXCHARDISPMODE1_IN                      : in   std_logic;
    TXCHARDISPVAL0_IN                       : in   std_logic;
    TXCHARDISPVAL1_IN                       : in   std_logic;
    TXCHARISK0_IN                           : in   std_logic;
    TXCHARISK1_IN                           : in   std_logic;
    ------------- Transmit Ports - TX Buffering and Phase Alignment ------------
    TXBUFSTATUS0_OUT                        : out  std_logic_vector(1 downto 0);
    TXBUFSTATUS1_OUT                        : out  std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TXDATA0_IN                              : in   std_logic_vector(7 downto 0);
    TXDATA1_IN                              : in   std_logic_vector(7 downto 0);
    TXOUTCLK0_OUT                           : out  std_logic;
    TXOUTCLK1_OUT                           : out  std_logic;
    TXRESET0_IN                             : in   std_logic;
    TXRESET1_IN                             : in   std_logic;
    TXUSRCLK0_IN                            : in   std_logic;
    TXUSRCLK1_IN                            : in   std_logic;
    TXUSRCLK20_IN                           : in   std_logic;
    TXUSRCLK21_IN                           : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TXN0_OUT                                : out  std_logic;
    TXN1_OUT                                : out  std_logic;
    TXP0_OUT                                : out  std_logic;
    TXP1_OUT                                : out  std_logic;
    -- Polarity control (DMN addition)
    rxpolarity: in std_logic_vector(1 downto 0);
    txpolarity: in std_logic_vector(1 downto 0)

);
end ROCKETIO_WRAPPER_GTX_TILE;

architecture RTL of ROCKETIO_WRAPPER_GTX_TILE is
    
--**************************** Signal Declarations ****************************

    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;

   

    -- RX Datapath signals
    signal rxdata0_i                        :   std_logic_vector(31 downto 0);
    signal rxchariscomma0_float_i           :   std_logic_vector(2 downto 0);
    signal rxcharisk0_float_i               :   std_logic_vector(2 downto 0);
    signal rxdisperr0_float_i               :   std_logic_vector(2 downto 0);
    signal rxnotintable0_float_i            :   std_logic_vector(2 downto 0);
    signal rxrundisp0_float_i               :   std_logic_vector(2 downto 0);

    -- TX Datapath signals
    signal txdata0_i                        :   std_logic_vector(31 downto 0);

   

    -- RX Datapath signals
    signal rxdata1_i                        :   std_logic_vector(31 downto 0);
    signal rxchariscomma1_float_i           :   std_logic_vector(2 downto 0);
    signal rxcharisk1_float_i               :   std_logic_vector(2 downto 0);
    signal rxdisperr1_float_i               :   std_logic_vector(2 downto 0);
    signal rxnotintable1_float_i            :   std_logic_vector(2 downto 0);
    signal rxrundisp1_float_i               :   std_logic_vector(2 downto 0);

    -- TX Datapath signals
    signal txdata1_i                        :   std_logic_vector(31 downto 0);




--******************************** Main Body of Code***************************
                       
begin                      

    ---------------------------  Static signal Assignments ---------------------   

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
     
    -------------------  GTP Datapath byte mapping  -----------------    

    RXDATA0_OUT    <=   rxdata0_i(7 downto 0);
    
    txdata0_i    <=   (tied_to_ground_vec_i(23 downto 0) & TXDATA0_IN);    

    RXDATA1_OUT    <=   rxdata1_i(7 downto 0);
    
    txdata1_i    <=   (tied_to_ground_vec_i(23 downto 0) & TXDATA1_IN);    




    ----------------------------- GTP_DUAL Instance  --------------------------   

    gtx_dual_i:GTX_DUAL
    generic map
    (

        --_______________________ Simulation-Only Attributes ___________________

        SIM_GTXRESET_SPEEDUP        =>       TILE_SIM_GTXRESET_SPEEDUP,
        SIM_PLL_PERDIV2             =>       TILE_SIM_PLL_PERDIV2,
        SIM_MODE                    =>       "FAST",
        SIM_RECEIVER_DETECT_PASS_0  =>       TRUE,
        SIM_RECEIVER_DETECT_PASS_1  =>       TRUE,

        --___________________________ Shared Attributes ________________________

        -------------------------- Tile and PLL Attributes ---------------------

        CLK25_DIVIDER               =>       5, 
        CLKINDC_B                   =>       TRUE,
        CLKRCV_TRST                 =>       TRUE,
        OOB_CLK_DIVIDER             =>       4,
        OVERSAMPLE_MODE             =>       FALSE,
        PLL_COM_CFG                 =>       x"21680a",
        PLL_CP_CFG                  =>       x"00",
        PLL_DIVSEL_FB               =>       4,
        PLL_DIVSEL_REF              =>       1,
        PLL_FB_DCCEN                =>       FALSE,
        PLL_LKDET_CFG               =>       "101",
        PLL_TDCC_CFG                =>       "000",
        PMA_COM_CFG                 =>       x"000000000000000000",


        --____________________ Transmit Interface Attributes ___________________


        ------------------- TX Buffering and Phase Alignment -------------------   

        TX_BUFFER_USE_0             =>       TRUE,
        TX_XCLK_SEL_0               =>       "TXOUT",
        TXRX_INVERT_0               =>       "011",        

        TX_BUFFER_USE_1             =>       TRUE,
        TX_XCLK_SEL_1               =>       "TXOUT",
        TXRX_INVERT_1               =>       "011",        

        --------------------- TX Gearbox Settings -----------------------------

        GEARBOX_ENDEC_0             =>       "000", 
        TXGEARBOX_USE_0            =>        FALSE,

        GEARBOX_ENDEC_1            =>        "000", 
        TXGEARBOX_USE_1            =>        FALSE,

        --------------------- TX Serial Line Rate settings ---------------------   

        PLL_TXDIVSEL_OUT_0          =>       4,

        PLL_TXDIVSEL_OUT_1          =>       4,

        --------------------- TX Driver and OOB signalling --------------------  

        CM_TRIM_0                   =>       "10",
        PMA_TX_CFG_0                =>       x"80082",
        TX_DETECT_RX_CFG_0          =>       x"1832",
        TX_IDLE_DELAY_0             =>       "010",

        CM_TRIM_1                   =>       "10",
        PMA_TX_CFG_1                =>       x"80082",
        TX_DETECT_RX_CFG_1          =>       x"1832",
        TX_IDLE_DELAY_1             =>       "010",

        ------------------ TX Pipe Control for PCI Express/SATA ---------------

        COM_BURST_VAL_0             =>       "1111",

        COM_BURST_VAL_1             =>       "1111",
        --_______________________ Receive Interface Attributes ________________


        ------------ RX Driver,OOB signalling,Coupling and Eq,CDR -------------  

        AC_CAP_DIS_0                =>       TRUE,
        OOBDETECT_THRESHOLD_0       =>       "111",
        PMA_CDR_SCAN_0              =>       x"6404035",
        PMA_RX_CFG_0                =>       x"0f44088",
        RCV_TERM_GND_0              =>       FALSE,
        RCV_TERM_VTTRX_0            =>       TRUE,
        TERMINATION_IMP_0           =>       50,

        AC_CAP_DIS_1                =>       TRUE,
        OOBDETECT_THRESHOLD_1       =>       "111",
        PMA_CDR_SCAN_1              =>       x"6404035",
        PMA_RX_CFG_1                =>       x"0f44088",  
        RCV_TERM_GND_1              =>       FALSE,
        RCV_TERM_VTTRX_1            =>       TRUE,
        TERMINATION_IMP_1           =>       50,

        TERMINATION_CTRL            =>       "10100",
        TERMINATION_OVRD            =>       FALSE,

        ---------------- RX Decision Feedback Equalizer(DFE)  ----------------  

        DFE_CFG_0                   =>       "1001111011",
                 
        DFE_CFG_1                   =>       "1001111011",

        DFE_CAL_TIME                =>       "00110",

        --------------------- RX Serial Line Rate Attributes ------------------   

        PLL_RXDIVSEL_OUT_0          =>       4,
        PLL_SATA_0                  =>       FALSE,

        PLL_RXDIVSEL_OUT_1          =>       4,
        PLL_SATA_1                  =>       FALSE,

        ----------------------- PRBS Detection Attributes ---------------------  

        PRBS_ERR_THRESHOLD_0        =>       x"00000001",

        PRBS_ERR_THRESHOLD_1        =>       x"00000001",

        ---------------- Comma Detection and Alignment Attributes -------------  

        ALIGN_COMMA_WORD_0          =>       1,
        COMMA_10B_ENABLE_0          =>       "0001111111",
        COMMA_DOUBLE_0              =>       FALSE,
        DEC_MCOMMA_DETECT_0         =>       TRUE,
        DEC_PCOMMA_DETECT_0         =>       TRUE,
        DEC_VALID_COMMA_ONLY_0      =>       FALSE,
        MCOMMA_10B_VALUE_0          =>       "1010000011",
        MCOMMA_DETECT_0             =>       TRUE,
        PCOMMA_10B_VALUE_0          =>       "0101111100",
        PCOMMA_DETECT_0             =>       TRUE,
        RX_SLIDE_MODE_0             =>       "PCS",

        ALIGN_COMMA_WORD_1          =>       1,
        COMMA_10B_ENABLE_1          =>       "0001111111",
        COMMA_DOUBLE_1              =>       FALSE,
        DEC_MCOMMA_DETECT_1         =>       TRUE,
        DEC_PCOMMA_DETECT_1         =>       TRUE,
        DEC_VALID_COMMA_ONLY_1      =>       FALSE,
        MCOMMA_10B_VALUE_1          =>       "1010000011",
        MCOMMA_DETECT_1             =>       TRUE,
        PCOMMA_10B_VALUE_1          =>       "0101111100",
        PCOMMA_DETECT_1             =>       TRUE,
        RX_SLIDE_MODE_1             =>       "PCS",

        ------------------ RX Loss-of-sync State Machine Attributes -----------  

        RX_LOSS_OF_SYNC_FSM_0       =>       FALSE,
        RX_LOS_INVALID_INCR_0       =>       8,
        RX_LOS_THRESHOLD_0          =>       128,

        RX_LOSS_OF_SYNC_FSM_1       =>       FALSE,
        RX_LOS_INVALID_INCR_1       =>       8,
        RX_LOS_THRESHOLD_1          =>       128,

        --------------------- RX Gearbox Settings -----------------------------

        RXGEARBOX_USE_0             =>       FALSE,

        RXGEARBOX_USE_1             =>       FALSE,

        -------------- RX Elastic Buffer and Phase alignment Attributes -------   

        PMA_RXSYNC_CFG_0            =>       x"00",
        RX_BUFFER_USE_0             =>       TRUE,
        RX_XCLK_SEL_0               =>       "RXREC",

        PMA_RXSYNC_CFG_1            =>       x"00",
        RX_BUFFER_USE_1             =>       TRUE,
        RX_XCLK_SEL_1               =>       "RXREC",                   

        ------------------------ Clock Correction Attributes ------------------   

        CLK_CORRECT_USE_0           =>       TRUE,
        CLK_COR_ADJ_LEN_0           =>       2,
        CLK_COR_DET_LEN_0           =>       2,
        CLK_COR_INSERT_IDLE_FLAG_0  =>       FALSE,
        CLK_COR_KEEP_IDLE_0         =>       FALSE,
        CLK_COR_MAX_LAT_0           =>       20,
        CLK_COR_MIN_LAT_0           =>       16,
        CLK_COR_PRECEDENCE_0        =>       TRUE,
        CLK_COR_REPEAT_WAIT_0       =>       0,
        CLK_COR_SEQ_1_1_0           =>       "0110111100",
        CLK_COR_SEQ_1_2_0           =>       "0001010000",
        CLK_COR_SEQ_1_3_0           =>       "0000000000",
        CLK_COR_SEQ_1_4_0           =>       "0000000000",
        CLK_COR_SEQ_1_ENABLE_0      =>       "0011",
        CLK_COR_SEQ_2_1_0           =>       "0110111100",
        CLK_COR_SEQ_2_2_0           =>       "0010110101",
        CLK_COR_SEQ_2_3_0           =>       "0000000000",
        CLK_COR_SEQ_2_4_0           =>       "0000000000",
        CLK_COR_SEQ_2_ENABLE_0      =>       "0011",
        CLK_COR_SEQ_2_USE_0         =>       TRUE,
        RX_DECODE_SEQ_MATCH_0       =>       TRUE,

        CLK_CORRECT_USE_1           =>       TRUE,
        CLK_COR_ADJ_LEN_1           =>       2,
        CLK_COR_DET_LEN_1           =>       2,
        CLK_COR_INSERT_IDLE_FLAG_1  =>       FALSE,
        CLK_COR_KEEP_IDLE_1         =>       FALSE,
        CLK_COR_MAX_LAT_1           =>       20,
        CLK_COR_MIN_LAT_1           =>       16,
        CLK_COR_PRECEDENCE_1        =>       TRUE,
        CLK_COR_REPEAT_WAIT_1       =>       0,
        CLK_COR_SEQ_1_1_1           =>       "0110111100",
        CLK_COR_SEQ_1_2_1           =>       "0001010000",
        CLK_COR_SEQ_1_3_1           =>       "0000000000",
        CLK_COR_SEQ_1_4_1           =>       "0000000000",
        CLK_COR_SEQ_1_ENABLE_1      =>       "0011",
        CLK_COR_SEQ_2_1_1           =>       "0110111100",
        CLK_COR_SEQ_2_2_1           =>       "0010110101",
        CLK_COR_SEQ_2_3_1           =>       "0000000000",
        CLK_COR_SEQ_2_4_1           =>       "0000000000",
        CLK_COR_SEQ_2_ENABLE_1      =>       "0011",
        CLK_COR_SEQ_2_USE_1         =>       TRUE,
        RX_DECODE_SEQ_MATCH_1       =>       TRUE,

        ------------------------ Channel Bonding Attributes -------------------   

        CB2_INH_CC_PERIOD_0         =>       8,
        CHAN_BOND_1_MAX_SKEW_0      =>       1,
        CHAN_BOND_2_MAX_SKEW_0      =>       1,
        CHAN_BOND_KEEP_ALIGN_0      =>       FALSE,
        CHAN_BOND_LEVEL_0           =>       TILE_CHAN_BOND_LEVEL_0,
        CHAN_BOND_MODE_0            =>       TILE_CHAN_BOND_MODE_0,
        CHAN_BOND_SEQ_1_1_0         =>       "0000000000",
        CHAN_BOND_SEQ_1_2_0         =>       "0000000000",
        CHAN_BOND_SEQ_1_3_0         =>       "0000000000",
        CHAN_BOND_SEQ_1_4_0         =>       "0000000000",
        CHAN_BOND_SEQ_1_ENABLE_0    =>       "0000",
        CHAN_BOND_SEQ_2_1_0         =>       "0000000000",
        CHAN_BOND_SEQ_2_2_0         =>       "0000000000",
        CHAN_BOND_SEQ_2_3_0         =>       "0000000000",
        CHAN_BOND_SEQ_2_4_0         =>       "0000000000",
        CHAN_BOND_SEQ_2_ENABLE_0    =>       "0000",
        CHAN_BOND_SEQ_2_USE_0       =>       FALSE,  
        CHAN_BOND_SEQ_LEN_0         =>       1,
        PCI_EXPRESS_MODE_0          =>       FALSE,   
     
        CB2_INH_CC_PERIOD_1         =>       8,
        CHAN_BOND_1_MAX_SKEW_1      =>       1,
        CHAN_BOND_2_MAX_SKEW_1      =>       1,
        CHAN_BOND_KEEP_ALIGN_1      =>       FALSE,
        CHAN_BOND_LEVEL_1           =>       TILE_CHAN_BOND_LEVEL_1,
        CHAN_BOND_MODE_1            =>       TILE_CHAN_BOND_MODE_1,
        CHAN_BOND_SEQ_1_1_1         =>       "0000000000",
        CHAN_BOND_SEQ_1_2_1         =>       "0000000000",
        CHAN_BOND_SEQ_1_3_1         =>       "0000000000",
        CHAN_BOND_SEQ_1_4_1         =>       "0000000000",
        CHAN_BOND_SEQ_1_ENABLE_1    =>       "0000",
        CHAN_BOND_SEQ_2_1_1         =>       "0000000000",
        CHAN_BOND_SEQ_2_2_1         =>       "0000000000",
        CHAN_BOND_SEQ_2_3_1         =>       "0000000000",
        CHAN_BOND_SEQ_2_4_1         =>       "0000000000",
        CHAN_BOND_SEQ_2_ENABLE_1    =>       "0000",
        CHAN_BOND_SEQ_2_USE_1       =>       FALSE,  
        CHAN_BOND_SEQ_LEN_1         =>       1,
        PCI_EXPRESS_MODE_1          =>       FALSE,

        -------- RX Attributes to Control Reset after Electrical Idle  ------

        RX_EN_IDLE_HOLD_DFE_0       =>       TRUE,
        RX_EN_IDLE_RESET_BUF_0      =>       TRUE,
        RX_IDLE_HI_CNT_0            =>       "1000",
        RX_IDLE_LO_CNT_0            =>       "0000",

        RX_EN_IDLE_HOLD_DFE_1       =>       TRUE,
        RX_EN_IDLE_RESET_BUF_1      =>       TRUE,
        RX_IDLE_HI_CNT_1            =>       "1000",
        RX_IDLE_LO_CNT_1            =>       "0000",


        CDR_PH_ADJ_TIME             =>       "01010",
        RX_EN_IDLE_RESET_FR         =>       TRUE,
        RX_EN_IDLE_HOLD_CDR         =>       FALSE,
        RX_EN_IDLE_RESET_PH         =>       TRUE,

        ------------------ RX Attributes for PCI Express/SATA ---------------

        RX_STATUS_FMT_0             =>       "PCIE",
        SATA_BURST_VAL_0            =>       "100",
        SATA_IDLE_VAL_0             =>       "100",
        SATA_MAX_BURST_0            =>       9,
        SATA_MAX_INIT_0             =>       27,
        SATA_MAX_WAKE_0             =>       9,
        SATA_MIN_BURST_0            =>       5,
        SATA_MIN_INIT_0             =>       15,
        SATA_MIN_WAKE_0             =>       5,
        TRANS_TIME_FROM_P2_0        =>       x"003c",
        TRANS_TIME_NON_P2_0         =>       x"0019",
        TRANS_TIME_TO_P2_0          =>       x"0064",

        RX_STATUS_FMT_1             =>       "PCIE",
        SATA_BURST_VAL_1            =>       "100",
        SATA_IDLE_VAL_1             =>       "100",
        SATA_MAX_BURST_1            =>       9,
        SATA_MAX_INIT_1             =>       27,
        SATA_MAX_WAKE_1             =>       9,
        SATA_MIN_BURST_1            =>       5,
        SATA_MIN_INIT_1             =>       15,
        SATA_MIN_WAKE_1             =>       5,
        TRANS_TIME_FROM_P2_1        =>       x"003c",
        TRANS_TIME_NON_P2_1         =>       x"0019",
        TRANS_TIME_TO_P2_1          =>       x"0064"
    ) 
    port map 
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK0                       =>      LOOPBACK0_IN,
        LOOPBACK1                       =>      LOOPBACK1_IN,

        RXPOWERDOWN0                    =>      RXPOWERDOWN0_IN,
        RXPOWERDOWN1                    =>      RXPOWERDOWN1_IN,
        TXPOWERDOWN0                    =>      TXPOWERDOWN0_IN,
        TXPOWERDOWN1                    =>      TXPOWERDOWN1_IN,       
        -------------- Receive Ports - 64b66b and 64b67b Gearbox Ports -------------
        RXDATAVALID0                    =>      open,
        RXDATAVALID1                    =>      open,
        RXGEARBOXSLIP0                  =>      tied_to_ground_i,
        RXGEARBOXSLIP1                  =>      tied_to_ground_i,
        RXHEADER0                       =>      open,
        RXHEADER1                       =>      open,
        RXHEADERVALID0                  =>      open,
        RXHEADERVALID1                  =>      open,
        RXSTARTOFSEQ0                   =>      open,
        RXSTARTOFSEQ1                   =>      open,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA0(3 downto 1)      =>      rxchariscomma0_float_i,
        RXCHARISCOMMA0(0)               =>      RXCHARISCOMMA0_OUT,
        RXCHARISK0(3 downto 1)          =>      rxcharisk0_float_i,
        RXCHARISK0(0)                   =>      RXCHARISK0_OUT,
        RXDEC8B10BUSE0                  =>      tied_to_vcc_i,
        RXDISPERR0(3 downto 1)          =>      rxdisperr0_float_i,
        RXDISPERR0(0)                   =>      RXDISPERR0_OUT,
        RXNOTINTABLE0(3 downto 1)       =>      rxnotintable0_float_i,
        RXNOTINTABLE0(0)                =>      RXNOTINTABLE0_OUT,
        RXRUNDISP0(3 downto 1)          =>      rxrundisp0_float_i,
        RXRUNDISP0(0)                   =>      RXRUNDISP0_OUT,
        RXCHARISCOMMA1(3 downto 1)      =>      rxchariscomma1_float_i,
        RXCHARISCOMMA1(0)               =>      RXCHARISCOMMA1_OUT,
        RXCHARISK1(3 downto 1)          =>      rxcharisk1_float_i,
        RXCHARISK1(0)                   =>      RXCHARISK1_OUT,
        RXDEC8B10BUSE1                  =>      tied_to_vcc_i,
        RXDISPERR1(3 downto 1)          =>      rxdisperr1_float_i,
        RXDISPERR1(0)                   =>      RXDISPERR1_OUT,
        RXNOTINTABLE1(3 downto 1)       =>      rxnotintable1_float_i,
        RXNOTINTABLE1(0)                =>      RXNOTINTABLE1_OUT,
        RXRUNDISP1(3 downto 1)          =>      rxrundisp1_float_i,
        RXRUNDISP1(0)                   =>      RXRUNDISP1_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ0                  =>      open,
        RXCHANBONDSEQ1                  =>      open,
        RXCHBONDI0                      =>      tied_to_ground_vec_i(3 downto 0),
        RXCHBONDI1                      =>      tied_to_ground_vec_i(3 downto 0),
        RXCHBONDO0                      =>      open,
        RXCHBONDO1                      =>      open,
        RXENCHANSYNC0                   =>      tied_to_ground_i,
        RXENCHANSYNC1                   =>      tied_to_ground_i,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT0                    =>      RXCLKCORCNT0_OUT,
        RXCLKCORCNT1                    =>      RXCLKCORCNT1_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED0                =>      open,
        RXBYTEISALIGNED1                =>      open,
        RXBYTEREALIGN0                  =>      open,
        RXBYTEREALIGN1                  =>      open,
        RXCOMMADET0                     =>      open,
        RXCOMMADET1                     =>      open,
        RXCOMMADETUSE0                  =>      tied_to_vcc_i,
        RXCOMMADETUSE1                  =>      tied_to_vcc_i,
        RXENMCOMMAALIGN0                =>      RXENMCOMMAALIGN0_IN,
        RXENMCOMMAALIGN1                =>      RXENMCOMMAALIGN1_IN,
        RXENPCOMMAALIGN0                =>      RXENPCOMMAALIGN0_IN,
        RXENPCOMMAALIGN1                =>      RXENPCOMMAALIGN1_IN,
        RXSLIDE0                        =>      tied_to_ground_i,
        RXSLIDE1                        =>      tied_to_ground_i,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        PRBSCNTRESET0                   =>      tied_to_ground_i,
        PRBSCNTRESET1                   =>      tied_to_ground_i,
        RXENPRBSTST0                    =>      tied_to_ground_vec_i(1 downto 0),
        RXENPRBSTST1                    =>      tied_to_ground_vec_i(1 downto 0),
        RXPRBSERR0                      =>      open,
        RXPRBSERR1                      =>      open,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA0                         =>      rxdata0_i,
        RXDATA1                         =>      rxdata1_i,
        RXDATAWIDTH0                    =>      "00",
        RXDATAWIDTH1                    =>      "00",
        RXRECCLK0                       =>      RXRECCLK0_OUT,
        RXRECCLK1                       =>      RXRECCLK1_OUT,
        RXRESET0                        =>      RXRESET0_IN,
        RXRESET1                        =>      RXRESET1_IN,
        RXUSRCLK0                       =>      RXUSRCLK0_IN,
        RXUSRCLK1                       =>      RXUSRCLK1_IN,
        RXUSRCLK20                      =>      RXUSRCLK20_IN,
        RXUSRCLK21                      =>      RXUSRCLK21_IN,
        ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
        DFECLKDLYADJ0                   =>      tied_to_ground_vec_i(5 downto 0),
        DFECLKDLYADJ1                   =>      tied_to_ground_vec_i(5 downto 0),
        DFECLKDLYADJMONITOR0            =>      open,
        DFECLKDLYADJMONITOR1            =>      open,
        DFEEYEDACMONITOR0               =>      open,
        DFEEYEDACMONITOR1               =>      open,
        DFESENSCAL0                     =>      open,
        DFESENSCAL1                     =>      open,
        DFETAP10                        =>      tied_to_ground_vec_i(4 downto 0),
        DFETAP11                        =>      tied_to_ground_vec_i(4 downto 0),
        DFETAP1MONITOR0                 =>      open,
        DFETAP1MONITOR1                 =>      open,
        DFETAP20                        =>      tied_to_ground_vec_i(4 downto 0),
        DFETAP21                        =>      tied_to_ground_vec_i(4 downto 0),
        DFETAP2MONITOR0                 =>      open,
        DFETAP2MONITOR1                 =>      open,
        DFETAP30                        =>      tied_to_ground_vec_i(3 downto 0),
        DFETAP31                        =>      tied_to_ground_vec_i(3 downto 0),
        DFETAP3MONITOR0                 =>      open,
        DFETAP3MONITOR1                 =>      open,
        DFETAP40                        =>      tied_to_ground_vec_i(3 downto 0),
        DFETAP41                        =>      tied_to_ground_vec_i(3 downto 0),
        DFETAP4MONITOR0                 =>      open,
        DFETAP4MONITOR1                 =>      open,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET0                     =>      tied_to_ground_i,
        RXCDRRESET1                     =>      tied_to_ground_i,
        RXELECIDLE0                     =>      RXELECIDLE0_OUT,
        RXELECIDLE1                     =>      RXELECIDLE1_OUT,
        RXENEQB0                        =>      tied_to_ground_i,
        RXENEQB1                        =>      tied_to_ground_i,
        RXEQMIX0                        =>      "11",
        RXEQMIX1                        =>      "11",
        RXEQPOLE0                       =>      tied_to_ground_vec_i(3 downto 0),
        RXEQPOLE1                       =>      tied_to_ground_vec_i(3 downto 0),
        RXN0                            =>      RXN0_IN,
        RXN1                            =>      RXN1_IN,
        RXP0                            =>      RXP0_IN,
        RXP1                            =>      RXP1_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET0                     =>      RXBUFRESET0_IN,
        RXBUFRESET1                     =>      RXBUFRESET1_IN,
        RXBUFSTATUS0                    =>      RXBUFSTATUS0_OUT,
        RXBUFSTATUS1                    =>      RXBUFSTATUS1_OUT,
        RXCHANISALIGNED0                =>      open,
        RXCHANISALIGNED1                =>      open,
        RXCHANREALIGN0                  =>      open,
        RXCHANREALIGN1                  =>      open,
        RXENPMAPHASEALIGN0              =>      tied_to_ground_i,
        RXENPMAPHASEALIGN1              =>      tied_to_ground_i,
        RXPMASETPHASE0                  =>      tied_to_ground_i,
        RXPMASETPHASE1                  =>      tied_to_ground_i,
        RXSTATUS0                       =>      open,
        RXSTATUS1                       =>      open,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC0                   =>      open,
        RXLOSSOFSYNC1                   =>      open,
        ---------------------- Receive Ports - RX Oversampling ---------------------
        RXENSAMPLEALIGN0                =>      tied_to_ground_i,
        RXENSAMPLEALIGN1                =>      tied_to_ground_i,
        RXOVERSAMPLEERR0                =>      open,
        RXOVERSAMPLEERR1                =>      open,
        -------------- Receive Ports - RX Pipe Control for PCI Express -------------
        PHYSTATUS0                      =>      open,
        PHYSTATUS1                      =>      open,
        RXVALID0                        =>      open,
        RXVALID1                        =>      open,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        RXPOLARITY0                     =>      rxpolarity(0),
        RXPOLARITY1                     =>      rxpolarity(1),
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR                           =>      tied_to_ground_vec_i(6 downto 0),
        DCLK                            =>      tied_to_ground_i,
        DEN                             =>      tied_to_ground_i,
        DI                              =>      tied_to_ground_vec_i(15 downto 0),
        DO                              =>      open,
        DRDY                            =>      open,
        DWE                             =>      tied_to_ground_i,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        CLKIN                           =>      CLKIN_IN,
        GTXRESET                        =>      GTXRESET_IN,
        GTXTEST                         =>      "10000000000000",
        INTDATAWIDTH                    =>      tied_to_vcc_i,
        PLLLKDET                        =>      PLLLKDET_OUT,
        PLLLKDETEN                      =>      tied_to_vcc_i,
        PLLPOWERDOWN                    =>      tied_to_ground_i,
        REFCLKOUT                       =>      REFCLKOUT_OUT,
        REFCLKPWRDNB                    =>      tied_to_vcc_i,
        RESETDONE0                      =>      RESETDONE0_OUT,
        RESETDONE1                      =>      RESETDONE1_OUT,
        -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
        TXGEARBOXREADY0                 =>      open,
        TXGEARBOXREADY1                 =>      open,
        TXHEADER0                       =>      tied_to_ground_vec_i(2 downto 0),
        TXHEADER1                       =>      tied_to_ground_vec_i(2 downto 0),
        TXSEQUENCE0                     =>      tied_to_ground_vec_i(6 downto 0),
        TXSEQUENCE1                     =>      tied_to_ground_vec_i(6 downto 0),
        TXSTARTSEQ0                     =>      tied_to_ground_i,
        TXSTARTSEQ1                     =>      tied_to_ground_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXBYPASS8B10B0                  =>      tied_to_ground_vec_i(3 downto 0),
        TXBYPASS8B10B1                  =>      tied_to_ground_vec_i(3 downto 0),
        TXCHARDISPMODE0(3 downto 1)     =>      tied_to_ground_vec_i(2 downto 0),
        TXCHARDISPMODE0(0)              =>      TXCHARDISPMODE0_IN,
        TXCHARDISPMODE1(3 downto 1)     =>      tied_to_ground_vec_i(2 downto 0),
        TXCHARDISPMODE1(0)              =>      TXCHARDISPMODE1_IN,
        TXCHARDISPVAL0(3 downto 1)      =>      tied_to_ground_vec_i(2 downto 0),
        TXCHARDISPVAL0(0)               =>      TXCHARDISPVAL0_IN,
        TXCHARDISPVAL1(3 downto 1)      =>      tied_to_ground_vec_i(2 downto 0),
        TXCHARDISPVAL1(0)               =>      TXCHARDISPVAL1_IN,
        TXCHARISK0(3 downto 1)          =>      tied_to_ground_vec_i(2 downto 0),
        TXCHARISK0(0)                   =>      TXCHARISK0_IN,
        TXCHARISK1(3 downto 1)          =>      tied_to_ground_vec_i(2 downto 0),
        TXCHARISK1(0)                   =>      TXCHARISK1_IN,
        TXENC8B10BUSE0                  =>      tied_to_vcc_i,
        TXENC8B10BUSE1                  =>      tied_to_vcc_i,
        TXKERR0                         =>      open,
        TXKERR1                         =>      open,
        TXRUNDISP0                      =>      open,
        TXRUNDISP1                      =>      open,
        ------------- Transmit Ports - TX Buffering and Phase Alignment ------------
        TXBUFSTATUS0                    =>      TXBUFSTATUS0_OUT,
        TXBUFSTATUS1                    =>      TXBUFSTATUS1_OUT,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA0                         =>      txdata0_i,
        TXDATA1                         =>      txdata1_i,
        TXDATAWIDTH0                    =>      "00",
        TXDATAWIDTH1                    =>      "00",
        TXOUTCLK0                       =>      TXOUTCLK0_OUT,
        TXOUTCLK1                       =>      TXOUTCLK1_OUT,
        TXRESET0                        =>      TXRESET0_IN,
        TXRESET1                        =>      TXRESET1_IN,
        TXUSRCLK0                       =>      TXUSRCLK0_IN,
        TXUSRCLK1                       =>      TXUSRCLK1_IN,
        TXUSRCLK20                      =>      TXUSRCLK20_IN,
        TXUSRCLK21                      =>      TXUSRCLK21_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXBUFDIFFCTRL0                  =>      "101",
        TXBUFDIFFCTRL1                  =>      "101",
        TXDIFFCTRL0                     =>      "000",
        TXDIFFCTRL1                     =>      "000",
        TXINHIBIT0                      =>      tied_to_ground_i,
        TXINHIBIT1                      =>      tied_to_ground_i,
        TXN0                            =>      TXN0_OUT,
        TXN1                            =>      TXN1_OUT,
        TXP0                            =>      TXP0_OUT,
        TXP1                            =>      TXP1_OUT,
        TXPREEMPHASIS0                  =>      "0000",
        TXPREEMPHASIS1                  =>      "0000",
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXENPMAPHASEALIGN0              =>      tied_to_ground_i,
        TXENPMAPHASEALIGN1              =>      tied_to_ground_i,
        TXPMASETPHASE0                  =>      tied_to_ground_i,
        TXPMASETPHASE1                  =>      tied_to_ground_i,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXENPRBSTST0                    =>      tied_to_ground_vec_i(1 downto 0),
        TXENPRBSTST1                    =>      tied_to_ground_vec_i(1 downto 0),
        -------------------- Transmit Ports - TX Polarity Control ------------------
        TXPOLARITY0                     =>      txpolarity(0),
        TXPOLARITY1                     =>      txpolarity(1),
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXDETECTRX0                     =>      tied_to_ground_i,
        TXDETECTRX1                     =>      tied_to_ground_i,
        TXELECIDLE0                     =>      tied_to_ground_i,
        TXELECIDLE1                     =>      tied_to_ground_i,
        --------------------- Transmit Ports - TX Ports for SATA -------------------
        TXCOMSTART0                     =>      tied_to_ground_i,
        TXCOMSTART1                     =>      tied_to_ground_i,
        TXCOMTYPE0                      =>      tied_to_ground_i,
        TXCOMTYPE1                      =>      tied_to_ground_i

    );

end RTL;
